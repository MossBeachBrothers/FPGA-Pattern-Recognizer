//process output image based on NN 
//alter color of output pixels based on classification results

module display_mux (); endmodule 


