//Top Module for NN 

module top_module (



); 

//NPU instance

//Control Instance



endmodule 